work.mem(main) :8: :8:
